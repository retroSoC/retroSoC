
`ifndef MDD_CONFIG_DEF_SVH
`define MDD_CONFIG_DEF_SVH

`define USER_MSTR_WIDTH 5
`define USER_SLAV_WIDTH 8
`define USER_GPIO_NUM   16

`endif