`timescale 1ns / 1ps

module retrosoc_top (
    input  clk_i,
    input  rst_n_i,
    input  uart0_rx_i,
    output uart0_tx_o,
    inout  gpio_io0,
    inout  gpio_io1,
    inout  gpio_io2,
    output psram_sck_o,
    output psram_nss0_o,
    inout  psram_dat0_io,
    inout  psram_dat1_io,
    inout  psram_dat2_io,
    inout  psram_dat3_io,
    output spisd_sck_o,
    output spisd_nss_o,
    output spisd_mosi_o,
    input  spisd_miso_i,
    output i2s_mclk_o,
    output i2s_sclk_o,
    output i2s_lrck_o,
    output i2s_dacdat_o,
    input  i2s_adcdat_i,
    inout  i2c_scl_io,
    inout  i2c_sda_io,
    output uart1_tx_o,
    input  uart1_rx_i,
    output pwm_0_o,
    input  ps2_clk_i,
    input  ps2_dat_i,
    output qspi_sck_o,
    output qspi_nss0_o,
    inout  qspi_dat0_io,
    output spfs_sck_o,
    output spfs_nss_o,
    output spfs_mosi_o,
    input  spfs_miso_i
);

  wire s_sys_clk;
  wire s_aud_clk;
  clk_wiz_0 u_clk_wiz_0 (
      .clk_in1 (clk_i),
      .clk_out1(s_sys_clk),
      .clk_out2(s_aud_clk)
  );

  retrosoc_asic u_retrosoc (
      .xi_i_pad             (s_sys_clk),
      .xo_o_pad             (),
      .extclk_i_pad         (s_sys_clk),
      .audclk_i_pad         (s_aud_clk),
      .irq_pin_i_pad        (1'b0),
`ifdef CORE_MDD
      .core_mdd_sel_0_i_pad (1'b0),
      .core_mdd_sel_1_i_pad (1'b0),
      .core_mdd_sel_2_i_pad (1'b0),
      .core_mdd_sel_3_i_pad (1'b0),
      .core_mdd_sel_4_i_pad (1'b0),
`endif
`ifdef IP_MDD
      .ip_mdd_gpio_0_io_pad (),
      .ip_mdd_gpio_1_io_pad (),
      .ip_mdd_gpio_2_io_pad (),
      .ip_mdd_gpio_3_io_pad (),
      .ip_mdd_gpio_4_io_pad (),
      .ip_mdd_gpio_5_io_pad (),
      .ip_mdd_gpio_6_io_pad (),
      .ip_mdd_gpio_7_io_pad (),
      .ip_mdd_gpio_8_io_pad (),
      .ip_mdd_gpio_9_io_pad (),
      .ip_mdd_gpio_10_io_pad(),
      .ip_mdd_gpio_11_io_pad(),
      .ip_mdd_gpio_12_io_pad(),
      .ip_mdd_gpio_13_io_pad(),
      .ip_mdd_gpio_14_io_pad(),
      .ip_mdd_gpio_15_io_pad(),
`endif
`ifdef HAVE_PLL
      .pll_cfg_0_i_pad      (1'b0),
      .pll_cfg_1_i_pad      (1'b0),
      .pll_cfg_2_i_pad      (1'b0),
`endif
      .clk_bypass_i_pad     (1'b1),
      .ext_rst_n_i_pad      (rst_n_i),
      .uart0_tx_o_pad       (uart0_tx_o),
      .uart0_rx_i_pad       (uart0_rx_i),
      .gpio_0_io_pad        (gpio_io0),
      .gpio_1_io_pad        (gpio_io1),
      .gpio_2_io_pad        (gpio_io2),
      .gpio_3_io_pad        (),
      .gpio_4_io_pad        (),
      .gpio_5_io_pad        (),
      .gpio_6_io_pad        (),
      .gpio_7_io_pad        (),
      .psram_sck_o_pad      (psram_sck_o),
      .psram_nss0_o_pad     (psram_nss0_o),
      .psram_nss1_o_pad     (),
      .psram_nss2_o_pad     (),
      .psram_nss3_o_pad     (),
      .psram_dat0_io_pad    (psram_dat0_io),
      .psram_dat1_io_pad    (psram_dat1_io),
      .psram_dat2_io_pad    (psram_dat2_io),
      .psram_dat3_io_pad    (psram_dat3_io),
      .spisd_sck_o_pad      (spisd_sck_o),
      .spisd_nss_o_pad      (spisd_nss_o),
      .spisd_mosi_o_pad     (spisd_mosi_o),
      .spisd_miso_i_pad     (spisd_miso_i),
      .i2s_mclk_o_pad       (),
      .i2s_sclk_o_pad       (),
      .i2s_lrck_o_pad       (),
      .i2s_dacdat_o_pad     (),
      .i2s_adcdat_i_pad     (),
      .uart1_tx_o_pad       (uart1_tx_o),
      .uart1_rx_i_pad       (uart1_rx_i),
      .pwm_0_o_pad          (pwm_0_o),
      .pwm_1_o_pad          (),
      .pwm_2_o_pad          (),
      .pwm_3_o_pad          (),
      .ps2_clk_i_pad        (ps2_clk_i),
      .ps2_dat_i_pad        (ps2_dat_i),
      .i2c_scl_io_pad       (i2c_scl_io),
      .i2c_sda_io_pad       (i2c_sda_io),
      .qspi_sck_o_pad       (qspi_sck_o),
      .qspi_nss0_o_pad      (qspi_nss0_o),
      .qspi_nss1_o_pad      (),
      .qspi_nss2_o_pad      (),
      .qspi_nss3_o_pad      (),
      .qspi_dat0_io_pad     (qspi_dat0_io),
      .qspi_dat1_io_pad     (),
      .qspi_dat2_io_pad     (),
      .qspi_dat3_io_pad     (),
      .spfs_sck_o_pad       (spfs_sck_o),
      .spfs_nss_o_pad       (spfs_nss_o),
      .spfs_mosi_o_pad      (spfs_mosi_o),
      .spfs_miso_i_pad      (spfs_miso_i)
  );
endmodule
