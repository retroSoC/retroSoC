// Copyright (c) 2023-2025 Yuchi Miao <miaoyuchi@ict.ac.cn>
// retroSoC is licensed under Mulan PSL v2.
// You can use this software according to the terms and conditions of the Mulan PSL v2.
// You may obtain a copy of Mulan PSL v2 at:
//             http://license.coscl.org.cn/MulanPSL2
// THIS SOFTWARE IS PROVIDED ON AN "AS IS" BASIS, WITHOUT WARRANTIES OF ANY KIND,
// EITHER EXPRESS OR IMPLIED, INCLUDING BUT NOT LIMITED TO NON-INFRINGEMENT,
// MERCHANTABILITY OR FIT FOR A PARTICULAR PURPOSE.
// See the Mulan PSL v2 for more details.


`include "mdd_config.svh"

module user_ip_wrapper (
    // verilog_format: off
    input  logic                        clk_i,
    input  logic                        rst_n_i,
    input  logic [`USER_SLAV_WIDTH-1:0] sel_i,
    user_gpio_if.dut                    gpio,
    apb4_if.slave                       apb
    // verilog_format: on
);

  // ====== GENERATED BY SCRIPT ======
  // verilog_format: off
  user_gpio_if u_user_1_gpio_if();
  user_gpio_if u_user_2_gpio_if();

  apb4_if u_user_1_apb_if(clk_i, rst_n_i);
  apb4_if u_user_2_apb_if(clk_i, rst_n_i);
  // ...
  // verilog_format: on
  always_comb begin
    gpio.gpio_out            = '0;
    gpio.gpio_oen            = '0;
    u_user_1_gpio_if.gpio_in = '0;
    u_user_2_gpio_if.gpio_in = '0;
    apb.pready               = '0;
    apb.prdata               = '0;
    u_user_1_apb_if.paddr    = '0;
    u_user_1_apb_if.pprot    = '0;
    u_user_1_apb_if.psel     = '0;
    u_user_1_apb_if.penable  = '0;
    u_user_1_apb_if.pwrite   = '0;
    u_user_1_apb_if.pwdata   = '0;
    u_user_1_apb_if.pstrb    = '0;
    u_user_2_apb_if.paddr    = '0;
    u_user_2_apb_if.pprot    = '0;
    u_user_2_apb_if.psel     = '0;
    u_user_2_apb_if.penable  = '0;
    u_user_2_apb_if.pwrite   = '0;
    u_user_2_apb_if.pwdata   = '0;
    u_user_2_apb_if.pstrb    = '0;
    unique case (sel_i)
      5'd1: begin
        gpio.gpio_out            = u_user_1_gpio_if.gpio_out;
        gpio.gpio_oen            = u_user_1_gpio_if.gpio_oen;
        u_user_1_gpio_if.gpio_in = gpio.gpio_in;
        apb.pready               = u_user_1_apb_if.pready;
        apb.prdata               = u_user_1_apb_if.prdata;
        u_user_1_apb_if.paddr    = apb.paddr;
        u_user_1_apb_if.pprot    = apb.pprot;
        u_user_1_apb_if.psel     = apb.psel;
        u_user_1_apb_if.penable  = apb.penable;
        u_user_1_apb_if.pwrite   = apb.pwrite;
        u_user_1_apb_if.pwdata   = apb.pwdata;
        u_user_1_apb_if.pstrb    = apb.pstrb;
      end
      5'd2: begin
        gpio.gpio_out            = u_user_2_gpio_if.gpio_out;
        gpio.gpio_oen            = u_user_2_gpio_if.gpio_oen;
        u_user_2_gpio_if.gpio_in = gpio.gpio_in;
        apb.pready               = u_user_2_apb_if.pready;
        apb.prdata               = u_user_2_apb_if.prdata;
        u_user_2_apb_if.paddr    = apb.paddr;
        u_user_2_apb_if.pprot    = apb.pprot;
        u_user_2_apb_if.psel     = apb.psel;
        u_user_2_apb_if.penable  = apb.penable;
        u_user_2_apb_if.pwrite   = apb.pwrite;
        u_user_2_apb_if.pwdata   = apb.pwdata;
        u_user_2_apb_if.pstrb    = apb.pstrb;
      end
      default: begin
        gpio.gpio_out            = '0;
        gpio.gpio_oen            = '0;
        u_user_1_gpio_if.gpio_in = '0;
        u_user_2_gpio_if.gpio_in = '0;
        apb.pready               = '0;
        apb.prdata               = '0;
        u_user_1_apb_if.paddr    = '0;
        u_user_1_apb_if.pprot    = '0;
        u_user_1_apb_if.psel     = '0;
        u_user_1_apb_if.penable  = '0;
        u_user_1_apb_if.pwrite   = '0;
        u_user_1_apb_if.pwdata   = '0;
        u_user_1_apb_if.pstrb    = '0;
        u_user_2_apb_if.paddr    = '0;
        u_user_2_apb_if.pprot    = '0;
        u_user_2_apb_if.psel     = '0;
        u_user_2_apb_if.penable  = '0;
        u_user_2_apb_if.pwrite   = '0;
        u_user_2_apb_if.pwdata   = '0;
        u_user_2_apb_if.pstrb    = '0;
      end
    endcase
  end

  user_ip_design #(1) u_user_1_ip_design (
      .clk_i  (clk_i),
      .rst_n_i(rst_n_i),
      .gpio   (u_user_1_gpio_if),
      .apb    (u_user_1_apb_if)
  );

  user_ip_design #(2) u_user_2_ip_design (
      .clk_i  (clk_i),
      .rst_n_i(rst_n_i),
      .gpio   (u_user_2_gpio_if),
      .apb    (u_user_2_apb_if)
  );

endmodule
